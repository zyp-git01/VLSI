module control (
    
);
    
endmodule