module output_select(
    input wire [3:0] select,
    
);












endmodule