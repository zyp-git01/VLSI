module compare #(
    parameter target_angle = 16'h500;
)
(
    input wire [15:0] 
);
    
endmodule